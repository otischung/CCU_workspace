//以前者(1ns)為單位，以後者(1ps)的時間，查看一次電路的行為
`timescale 1ns/1ps

//宣告module名稱,輸出入名稱
module lab9_optimized_serial_multiplier(
	clk, 
	rst, 
	in_a, 
	in_b, 
	Product, 
	Product_Valid
);
// in_a * in_b = Product
// in_a is Multiplicand , in_b is Multiplier
					
//定義port, 包含input, output
input clk, rst;
input [7:0] in_a;			// Multiplicand
input [7:0] in_b;			// Multiplier
output [15:0] Product;
output Product_Valid;

reg [7:0] Mplicand;		//被乘數
reg [7:0] Mplier;			//乘數
reg [15:0] Product;
reg Product_Valid;
reg [5:0] Counter;
reg sign;			//正負號判斷 (signed)

//Counter
always @(posedge clk or posedge rst) begin
	if (rst)
		Counter <= 6'b0;
	else
		Counter <= Counter + 6'b1;
end

//Product
always @(posedge clk or posedge rst) begin
	//初始化數值
	if (rst) begin
		Product <= 16'b0;
		Mplicand <= 16'b0;
		Mplier <= 8'b0;		
	end 
	//輸入乘數與被乘數
	else if (Counter == 6'd0) begin
		Mplicand <= in_a;
		Mplier <= in_b;
        Product <= { 8'b0, in_b };
	end 
	//乘法與數值移位
	else if (Counter <= 6'd8) begin
		if (Product[0] == 1'b1) begin  // LSB
            Product = Product + { Mplicand, 8'b0 };
        end
		Product = Product >> 1'b1;
	end 
	else begin
		Product <= Product;
		Mplicand <= Mplicand;
		Mplier <= Mplier;
	end
end

//Product_Valid
always @(posedge clk or posedge rst) begin
	if (rst)
		Product_Valid <=1'b0;
	else if (Counter == 6'd9)
		Product_Valid <=1'b1;
	else
		Product_Valid <=1'b0;
end

endmodule
